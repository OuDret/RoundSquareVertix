RECT -15.0 -25.0 15.0 25.0 ;
RECT -25.0 -15.0 -15.0 15.0 ;
RECT 15.0 -15.0 25.0 15.0 ;
RECT -15.5 15.0 -15.0 25.0 ;
RECT -15.5 -25.0 -15.0 -15.0 ;
RECT 15.0 15.0 15.5 25.0 ;
RECT 15.0 -25.0 15.5 -15.0 ;
RECT -16.0 15.0 -15.5 24.99 ;
RECT -16.0 -24.99 -15.5 -15.0 ;
RECT 15.5 15.0 16.0 24.99 ;
RECT 15.5 -24.99 16.0 -15.0 ;
RECT -16.5 15.0 -16.0 24.95 ;
RECT -16.5 -24.95 -16.0 -15.0 ;
RECT 16.0 15.0 16.5 24.95 ;
RECT 16.0 -24.95 16.5 -15.0 ;
RECT -17.0 15.0 -16.5 24.89 ;
RECT -17.0 -24.89 -16.5 -15.0 ;
RECT 16.5 15.0 17.0 24.89 ;
RECT 16.5 -24.89 17.0 -15.0 ;
RECT -17.5 15.0 -17.0 24.8 ;
RECT -17.5 -24.8 -17.0 -15.0 ;
RECT 17.0 15.0 17.5 24.8 ;
RECT 17.0 -24.8 17.5 -15.0 ;
RECT -18.0 15.0 -17.5 24.68 ;
RECT -18.0 -24.68 -17.5 -15.0 ;
RECT 17.5 15.0 18.0 24.68 ;
RECT 17.5 -24.68 18.0 -15.0 ;
RECT -18.5 15.0 -18.0 24.54 ;
RECT -18.5 -24.54 -18.0 -15.0 ;
RECT 18.0 15.0 18.5 24.54 ;
RECT 18.0 -24.54 18.5 -15.0 ;
RECT -19.0 15.0 -18.5 24.37 ;
RECT -19.0 -24.37 -18.5 -15.0 ;
RECT 18.5 15.0 19.0 24.37 ;
RECT 18.5 -24.37 19.0 -15.0 ;
RECT -19.5 15.0 -19.0 24.17 ;
RECT -19.5 -24.17 -19.0 -15.0 ;
RECT 19.0 15.0 19.5 24.17 ;
RECT 19.0 -24.17 19.5 -15.0 ;
RECT -20.0 15.0 -19.5 23.93 ;
RECT -20.0 -23.93 -19.5 -15.0 ;
RECT 19.5 15.0 20.0 23.93 ;
RECT 19.5 -23.93 20.0 -15.0 ;
RECT -20.5 15.0 -20.0 23.66 ;
RECT -20.5 -23.66 -20.0 -15.0 ;
RECT 20.0 15.0 20.5 23.66 ;
RECT 20.0 -23.66 20.5 -15.0 ;
RECT -21.0 15.0 -20.5 23.35 ;
RECT -21.0 -23.35 -20.5 -15.0 ;
RECT 20.5 15.0 21.0 23.35 ;
RECT 20.5 -23.35 21.0 -15.0 ;
RECT -21.5 15.0 -21.0 23.0 ;
RECT -21.5 -23.0 -21.0 -15.0 ;
RECT 21.0 15.0 21.5 23.0 ;
RECT 21.0 -23.0 21.5 -15.0 ;
RECT -22.0 15.0 -21.5 22.6 ;
RECT -22.0 -22.6 -21.5 -15.0 ;
RECT 21.5 15.0 22.0 22.6 ;
RECT 21.5 -22.6 22.0 -15.0 ;
RECT -22.5 15.0 -22.0 22.14 ;
RECT -22.5 -22.14 -22.0 -15.0 ;
RECT 22.0 15.0 22.5 22.14 ;
RECT 22.0 -22.14 22.5 -15.0 ;
RECT -23.0 15.0 -22.5 21.61 ;
RECT -23.0 -21.61 -22.5 -15.0 ;
RECT 22.5 15.0 23.0 21.61 ;
RECT 22.5 -21.61 23.0 -15.0 ;
RECT -23.5 15.0 -23.0 21.0 ;
RECT -23.5 -21.0 -23.0 -15.0 ;
RECT 23.0 15.0 23.5 21.0 ;
RECT 23.0 -21.0 23.5 -15.0 ;
RECT -24.0 15.0 -23.5 20.27 ;
RECT -24.0 -20.27 -23.5 -15.0 ;
RECT 23.5 15.0 24.0 20.27 ;
RECT 23.5 -20.27 24.0 -15.0 ;
RECT -24.5 15.0 -24.0 19.36 ;
RECT -24.5 -19.36 -24.0 -15.0 ;
RECT 24.0 15.0 24.5 19.36 ;
RECT 24.0 -19.36 24.5 -15.0 ;
RECT -25.0 15.0 -24.5 18.12 ;
RECT -25.0 -18.12 -24.5 -15.0 ;
RECT 24.5 15.0 25.0 18.12 ;
RECT 24.5 -18.12 25.0 -15.0 ;
